`include "mycpu.svh"

import mycpu_pkg::*;

module ir
  (
   input logic 	       clk,
   input logic 	       rst_n,
   input logic 	       il_in,
   input logic [15:0]  ins_in,
   output logic [15:0] ins_out,
   output logic [15:0] ia_out,
   output logic [15:0] iv_out   
   );
   
   
endmodule


